magic
tech sky130A
magscale 1 2
timestamp 1665597733
<< locali >>
rect 334 -166 528 -142
rect -44 -180 20 -166
rect -44 -214 -28 -180
rect 6 -214 20 -180
rect -44 -228 20 -214
rect 334 -322 362 -166
rect 502 -322 528 -166
rect 334 -344 528 -322
<< viali >>
rect -28 -214 6 -180
rect 362 -322 502 -166
rect 900 -224 968 -156
<< metal1 >>
rect 334 -166 528 -142
rect 894 -156 974 -150
rect -44 -180 20 -166
rect -44 -214 -28 -180
rect 6 -214 20 -180
rect -44 -228 20 -214
rect 334 -322 362 -166
rect 502 -322 528 -166
rect 888 -224 900 -156
rect 968 -224 980 -156
rect 894 -230 974 -224
rect 334 -344 528 -322
rect 1278 -543 1598 -164
rect 1278 -613 1757 -543
rect 1827 -613 1833 -543
rect 1278 -860 1598 -613
rect 1278 -1186 1598 -1180
<< via1 >>
rect 1757 -613 1827 -543
rect 1278 -1180 1598 -860
<< metal2 >>
rect 1757 -543 1827 -537
rect 1827 -613 1975 -543
rect 2045 -613 2054 -543
rect 1757 -619 1827 -613
rect 2663 -860 2973 -856
rect 1272 -1180 1278 -860
rect 1598 -865 2978 -860
rect 1598 -1175 2663 -865
rect 2973 -1175 2978 -865
rect 1598 -1180 2978 -1175
rect 2663 -1184 2973 -1180
<< via2 >>
rect 1975 -613 2045 -543
rect 2663 -1175 2973 -865
<< metal3 >>
rect 1975 -237 2045 -231
rect 1975 -538 2045 -307
rect 1970 -543 2050 -538
rect 1970 -613 1975 -543
rect 2045 -613 2050 -543
rect 1970 -618 2050 -613
rect 3757 -860 4075 -855
rect 2658 -861 4076 -860
rect 2658 -865 3757 -861
rect 2658 -1175 2663 -865
rect 2973 -1175 3757 -865
rect 2658 -1179 3757 -1175
rect 4075 -1179 4076 -861
rect 2658 -1180 4076 -1179
rect 3757 -1185 4075 -1180
<< via3 >>
rect 1975 -307 2045 -237
rect 3757 -1179 4075 -861
<< metal4 >>
rect 1974 -237 2046 -236
rect 1974 -307 1975 -237
rect 2045 -307 2392 -237
rect 1974 -308 2046 -307
rect 3756 -136 4076 -112
rect 3756 -408 3780 -136
rect 4052 -408 4076 -136
rect 3756 -861 4076 -408
rect 3756 -1179 3757 -861
rect 4075 -1179 4076 -861
rect 3756 -1180 4076 -1179
<< via4 >>
rect 2392 -432 2712 -112
rect 3780 -408 4052 -136
<< metal5 >>
rect 2368 -112 2736 -88
rect 2368 -432 2392 -112
rect 2712 -136 4076 -112
rect 2712 -408 3780 -136
rect 4052 -408 4076 -136
rect 2712 -432 4076 -408
rect 2368 -456 2736 -432
<< labels >>
flabel space -32 16 -32 16 0 FreeSans 320 0 0 0 Exercise_2a
flabel space -14 -74 -14 -74 0 FreeSans 320 0 0 0 Via_size
flabel space 440 14 440 14 0 FreeSans 320 0 0 0 Exercise_2b
flabel space 438 -66 438 -66 0 FreeSans 320 0 0 0 Multiple_vias
flabel space 948 4 948 4 0 FreeSans 320 0 0 0 Exercise_2c
flabel space 938 -68 938 -68 0 FreeSans 320 0 0 0 Via_overlap
flabel space 1540 -4 1540 -4 0 FreeSans 320 0 0 0 Exercise_2d
flabel space 1534 -66 1534 -66 0 FreeSans 320 0 0 0 Auto_generate_via
<< end >>
