magic
tech sky130A
magscale 1 2
timestamp 1665496688
<< metal1 >>
rect 922 1376 1122 1520
rect 730 1154 1366 1376
rect 730 1152 1278 1154
rect 672 1040 1040 1092
rect 672 788 724 1040
rect 1338 1008 1366 1154
rect 838 978 1366 1008
rect 1126 880 1166 888
rect 932 837 978 874
rect 1124 837 1170 880
rect 932 792 1309 837
rect 618 762 724 788
rect 618 720 1130 762
rect 618 686 680 720
rect 434 668 680 686
rect 322 646 680 668
rect 322 468 666 646
rect 504 466 666 468
rect 1264 554 1309 792
rect 1542 554 1742 700
rect 1264 510 1742 554
rect 614 286 664 466
rect 614 228 1040 286
rect 614 -38 664 228
rect 1264 199 1309 510
rect 1542 500 1742 510
rect 842 154 1309 199
rect 942 38 988 94
rect 1134 38 1180 96
rect 1238 38 1284 74
rect 936 -6 1284 38
rect 614 -72 1136 -38
rect 614 -74 664 -72
rect 876 -74 1136 -72
rect 1238 -136 1284 -6
rect 662 -176 1284 -136
rect 662 -286 1280 -176
rect 996 -472 1196 -286
use sky130_fd_pr__pfet_01v8_72SH2U  XM2
timestamp 1665427272
transform 1 0 1003 0 1 903
box -311 -319 311 319
use sky130_fd_pr__nfet_01v8_385SSZ  sky130_fd_pr__nfet_01v8_385SSZ_0
timestamp 1665427272
transform 1 0 1013 0 1 96
box -311 -310 311 310
<< labels >>
flabel metal1 922 1320 1122 1520 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 996 -472 1196 -272 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 322 468 522 668 0 FreeSans 256 0 0 0 in
port 2 nsew
flabel metal1 1542 500 1742 700 0 FreeSans 256 0 0 0 out
port 3 nsew
<< end >>
