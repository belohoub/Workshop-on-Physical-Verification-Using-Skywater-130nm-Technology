magic
tech sky130A
magscale 1 2
timestamp 1665496708
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -125 -147 -67 -141
rect 67 -147 125 -141
rect -125 -181 -113 -147
rect 67 -181 79 -147
rect -125 -187 -67 -181
rect 67 -187 125 -181
<< nwell >>
rect -311 -319 311 319
<< pmos >>
rect -114 -100 -78 100
rect -18 -100 18 100
rect 78 -100 114 100
<< pdiff >>
rect -173 88 -114 100
rect -173 -88 -161 88
rect -127 -88 -114 88
rect -173 -100 -114 -88
rect -78 88 -18 100
rect -78 -88 -65 88
rect -31 -88 -18 88
rect -78 -100 -18 -88
rect 18 88 78 100
rect 18 -88 31 88
rect 65 -88 78 88
rect 18 -100 78 -88
rect 114 88 173 100
rect 114 -88 127 88
rect 161 -88 173 88
rect 114 -100 173 -88
<< pdiffc >>
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
<< nsubdiff >>
rect -275 249 -179 283
rect 179 249 275 283
rect -275 187 -241 249
rect 241 187 275 249
rect -275 -249 -241 -187
rect 241 -249 275 -187
rect -275 -283 -179 -249
rect 179 -283 275 -249
<< nsubdiffcont >>
rect -179 249 179 283
rect -275 -187 -241 187
rect 241 -187 275 187
rect -179 -283 179 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -114 100 -78 126
rect -18 100 18 131
rect 78 100 114 126
rect -114 -131 -78 -100
rect -18 -126 18 -100
rect 78 -131 114 -100
rect -129 -147 -63 -131
rect -129 -181 -113 -147
rect -79 -181 -63 -147
rect -129 -197 -63 -181
rect 63 -147 129 -131
rect 63 -181 79 -147
rect 113 -181 129 -147
rect 63 -197 129 -181
<< polycont >>
rect -17 147 17 181
rect -113 -181 -79 -147
rect 79 -181 113 -147
<< locali >>
rect -275 249 -179 283
rect 179 249 275 283
rect -275 187 -241 249
rect 241 187 275 249
rect -33 147 -17 181
rect 17 147 33 181
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect -129 -181 -113 -147
rect -79 -181 -63 -147
rect 63 -181 79 -147
rect 113 -181 129 -147
rect -275 -249 -241 -187
rect 241 -249 275 -187
rect -275 -283 -179 -249
rect 179 -283 275 -249
<< viali >>
rect -17 147 17 181
rect -161 18 -127 71
rect -65 -26 -31 26
rect 31 18 65 71
rect 127 -26 161 26
rect -113 -181 -79 -147
rect 79 -181 113 -147
<< metal1 >>
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -167 71 -121 83
rect -167 18 -161 71
rect -127 18 -121 71
rect 25 71 71 83
rect -167 6 -121 18
rect -71 26 -25 38
rect -71 -26 -65 26
rect -31 -26 -25 26
rect 25 18 31 71
rect 65 18 71 71
rect 25 6 71 18
rect 121 26 167 38
rect -71 -38 -25 -26
rect 121 -26 127 26
rect 161 -26 167 26
rect 121 -38 167 -26
rect -125 -147 -67 -141
rect -125 -181 -113 -147
rect -79 -181 -67 -147
rect -125 -187 -67 -181
rect 67 -147 125 -141
rect 67 -181 79 -147
rect 113 -181 125 -147
rect 67 -187 125 -181
<< labels >>
rlabel pmos 17 9 17 9 1 S$
rlabel pmos -113 -3 -113 -3 1 S$
rlabel pmos 79 7 79 7 1 S$
<< properties >>
string FIXED_BBOX -258 -266 258 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.18 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn -30 viasrc 30
<< end >>
