magic
tech sky130A
magscale 1 2
timestamp 1665600495
<< dnwell >>
rect 2062 -1012 3088 -158
rect 2084 -1096 3088 -1012
rect 2084 -1100 3058 -1096
rect 4944 -1784 8098 1338
<< nwell >>
rect 4864 1132 8178 1418
rect -276 -476 -26 -184
rect 640 -436 890 -178
rect 1703 -365 3371 55
rect 1703 -806 2271 -365
rect 2877 -806 3371 -365
rect 1703 -890 3371 -806
rect 1700 -1370 3371 -890
rect 1700 -1374 3169 -1370
rect 4864 -1578 5150 1132
rect 7892 -1578 8178 1132
rect 4864 -1864 8178 -1578
<< pwell >>
rect 44 -434 294 -176
rect 960 -428 1210 -170
<< psubdiff >>
rect 1112 -222 1172 -192
rect 1112 -386 1118 -222
rect 1164 -386 1172 -222
rect 1112 -414 1172 -386
<< nsubdiff >>
rect 4901 1361 8141 1381
rect 4901 1327 4981 1361
rect 8061 1327 8141 1361
rect 4901 1307 8141 1327
rect 4901 1301 4975 1307
rect 682 -244 752 -214
rect -208 -290 -122 -264
rect -208 -402 -192 -290
rect -134 -402 -122 -290
rect 682 -374 698 -244
rect 738 -374 752 -244
rect 682 -400 752 -374
rect -208 -428 -122 -402
rect 2072 -1042 2352 -1020
rect 2072 -1084 2110 -1042
rect 2286 -1084 2352 -1042
rect 2072 -1106 2352 -1084
rect 4901 -1747 4921 1301
rect 4955 -1747 4975 1301
rect 4901 -1753 4975 -1747
rect 8067 1301 8141 1307
rect 8067 -1747 8087 1301
rect 8121 -1747 8141 1301
rect 8067 -1753 8141 -1747
rect 4901 -1773 8141 -1753
rect 4901 -1807 4981 -1773
rect 8061 -1807 8141 -1773
rect 4901 -1827 8141 -1807
<< psubdiffcont >>
rect 1118 -386 1164 -222
<< nsubdiffcont >>
rect 4981 1327 8061 1361
rect -192 -402 -134 -290
rect 698 -374 738 -244
rect 2110 -1084 2286 -1042
rect 4921 -1747 4955 1301
rect 8087 -1747 8121 1301
rect 4981 -1807 8061 -1773
<< locali >>
rect 4921 1327 4981 1361
rect 8061 1327 8121 1361
rect 4921 1301 4955 1327
rect 682 -244 752 -214
rect -192 -290 -134 -274
rect 682 -374 698 -244
rect 738 -374 752 -244
rect 682 -400 752 -374
rect 1118 -222 1164 -206
rect 1118 -402 1164 -386
rect -192 -418 -134 -402
rect 2086 -1084 2110 -1042
rect 2286 -1084 2310 -1042
rect 4921 -1773 4955 -1747
rect 8087 1301 8121 1327
rect 8087 -1773 8121 -1747
rect 4921 -1807 4981 -1773
rect 8061 -1807 8121 -1773
<< labels >>
flabel space -28 8 -28 8 0 FreeSans 320 0 0 0 Exercise_4a
flabel space -26 -68 -26 -68 0 FreeSans 320 0 0 0 Wells
flabel space 926 -16 926 -16 0 FreeSans 320 0 0 0 Exercise_4b
flabel space 920 -84 920 -84 0 FreeSans 320 0 0 0 Wells
flabel space 2158 196 2158 196 0 FreeSans 320 0 0 0 Exercise_4c
flabel space 2144 120 2144 120 0 FreeSans 320 0 0 0 Deep_NWell
<< end >>
