magic
tech sky130A
magscale 1 2
timestamp 1665598441
<< locali >>
rect -347 673 -108 707
rect -142 452 -108 673
<< viali >>
rect -381 673 -347 707
<< metal1 >>
rect -387 716 -341 719
rect -396 664 -390 716
rect -338 664 -332 716
rect -387 661 -341 664
rect 882 614 1192 698
rect 882 530 996 614
rect 1078 530 1192 614
rect 882 442 1192 530
<< via1 >>
rect -390 707 -338 716
rect -390 673 -381 707
rect -381 673 -347 707
rect -347 673 -338 707
rect -390 664 -338 673
<< metal2 >>
rect -664 901 -347 934
rect -380 716 -347 901
rect -396 664 -390 716
rect -338 664 -332 716
<< metal4 >>
rect 16 590 114 688
<< labels >>
flabel space 70 912 70 912 0 FreeSans 320 0 0 0 Exercise_3a
flabel space 64 828 64 828 0 FreeSans 320 0 0 0 Minimum_area_rule
flabel space 1042 944 1042 944 0 FreeSans 320 0 0 0 Exercise_3b
flabel space 1018 844 1018 844 0 FreeSans 320 0 0 0 Minimum_hole_rule
flabel space 1000 334 1000 334 0 FreeSans 320 0 0 0 *must_use_drc_style_sky130(full)*
<< end >>
