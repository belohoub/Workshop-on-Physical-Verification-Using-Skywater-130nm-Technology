* NGSPICE file created from all.ext - technology: sky130A

.subckt all vdd vss in out
X0 vdd in out XM2/w_n311_n319# sky130_fd_pr__pfet_01v8 ad=5.95e+11p pd=5.19e+06u as=5.95e+11p ps=5.19e+06u w=1e+06u l=180000u
X1 out in vdd XM2/w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X2 out in vdd XM2/w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X3 vss in out VSUBS sky130_fd_pr__nfet_01v8 ad=5.95e+11p pd=5.19e+06u as=5.95e+11p ps=5.19e+06u w=1e+06u l=180000u
X4 vss in out VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X5 out in vss VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends
