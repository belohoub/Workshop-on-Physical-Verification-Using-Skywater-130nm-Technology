magic
tech sky130A
magscale 1 2
timestamp 1665685298
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 -177 0 1 -1239
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  sky130_fd_sc_hd__nor2_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 -637 0 1 -1239
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 910 0 1 -1240
box -38 -48 130 592
<< labels >>
flabel space 88 -427 88 -427 0 FreeSans 320 0 0 0 Exercise_9a
flabel space 99 -494 99 -494 0 FreeSans 320 0 0 0 Latchup_rules
<< end >>
